`include "config.vh"

module overlay(
    input wire clk,
    input wire rst,
    input wire clk_2x,

    // inputs from controller
    input wire `Packet 

);
